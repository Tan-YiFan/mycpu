package forward_pkg;
    import common::*;
    typedef enum logic [1:0] {
        NOFORWARD,
        FORWARDM,
        FORWARDW
    } forward_t;
    
endpackage