//  Package: fetch_pkg
//
package fetch_pkg;
    //  Group: Typedefs
    typedef struct packed {
        word_t pcplus4;
        logic in_delay_slot;
    } fetch_data_t;
    

    //  Group: Parameters
    

    
endpackage: fetch_pkg
